module And (input wire branch, input wire zero, output wire saiAnd);

	assign saiAnd = branch & zero;
	
endmodule
